module alu_1bit (ctrl, busA, busB, zero, overflow, cout, cin, negative, out);
	input  logic [2:0]  ctrl;
	input  logic busA, busB;
	
   output logic out, negative, zero, overflow, cout;
	
	always_comb begin

	end

endmodule 